\m5_TLV_version 1d: tl-x.org
\m5
   
   // =================================================
   // Welcome!  New to Makerchip? Try the "Learn" menu.
   // =================================================
   
   //use(m5-1.0)   /// uncomment to use M5 macro library.
\SV
   // Macro providing required top-level module definition, random
   // stimulus support, and Verilator config.
   m5_makerchip_module   // (Expanded in Nav-TLV pane.)
\TLV
   $reset = *reset;
   
   $inv = ! $in1;
   $and = $in1 && $in2;
   $or = $in1 || $in2;
   $exor = $in1 ^ $in2 ;
   $nand = !( $in1 && $in2);
   $nor = !($in1 || $in2);
   $exnor = ! ($in1 ^ $in2) ;
   
   // Assert these to end simulation (before Makerchip cycle limit).
   *passed = *cyc_cnt > 40;
   *failed = 1'b0;
\SV
   endmodule
